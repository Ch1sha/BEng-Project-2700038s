/* verilator lint_off WIDTHEXPAND */
/* verilator lint_off BLKSEQ */
/* verilator lint_off REALCVT */
`define SINE_SIZE 8
`define TABLE_SIZE 32
`define TABLE_REG_SIZE 6
`define PHASE_SIZE 8 // resolution for phase input (from -180º to 180º)

module sine_wave (
    input logic clock, 
    input logic reset,
    input logic signed [`PHASE_SIZE:0] phase, // phase input determines the starting point of the sine wave, no -1 to handle signed values
    output logic [`SINE_SIZE-1:0] sine, // n-bit Sine wave output
    output integer phaseIdxOut,
    output integer i
);

    logic [`SINE_SIZE-1:0] sine_wave_table [0:`TABLE_SIZE-1]; // 50 samples of sine wave
    logic [`TABLE_REG_SIZE-1:0] logic_table_size;
    half_sine_table sine_table_inst (
        .sine_wave(sine_wave_table),
        .table_size(logic_table_size)
    );

    // Signal to hold the previous value of phase
    logic signed [`PHASE_SIZE:0] prev_phase;
    integer phaseIdx;
    integer tableSize;
    //integer i = phase; // Start from the given phase
    logic reverseTraversal = 0; // Reverse traversal flag

    // Function to calculate the starting index based on phase
    function integer calculate_start_index(input integer phaseIndex);
        integer midpoint;
        integer start_index;
        begin
            midpoint = (`TABLE_SIZE / 2); // Exact midpoint index of the sine table

            // Offset from midpoint
            start_index = midpoint + phaseIndex;

            // Ensure the index is positive
            if (start_index < 0) begin
                start_index = -start_index;
            end

            calculate_start_index = start_index;
        end
    endfunction

    // Takes in phase value in degrees and returns the corresponding phase value index for sine wave table
    function signed [`PHASE_SIZE:0] phase_to_phaseVal(input signed [`PHASE_SIZE:0] phaseIn);
        logic signed [`PHASE_SIZE:0] minVal; // Minimum phase value
        logic signed [`PHASE_SIZE:0] maxVal; // Maximum phase value = midpoint
        begin
            minVal = -3*(`TABLE_SIZE/2)+1;
            maxVal = (`TABLE_SIZE/2) -1;

            if (phaseIn >= 0 && phaseIn <= 90) begin
                // Map [0º, 90º] to [0, maxVal]
                phase_to_phaseVal = $floor(phaseIn * maxVal / 90);
            end
            else if (phaseIn > 90 && phaseIn <= 180) begin
                // Map [90º, 180º] to [minVal, -TABLE_SIZE]
                phase_to_phaseVal = minVal + $floor((phaseIn - 90) * maxVal / 90);
            end
            else if (phaseIn >= -180 && phaseIn < 0) begin
                // Map [-180º, 0º] to [TABLE_SIZE, 0]
                phase_to_phaseVal = -`TABLE_SIZE + $floor((phaseIn + 180) * `TABLE_SIZE / 180);
            end
            else begin
                // Clamp phase to valid range [-180º, 180º]
                phase_to_phaseVal = (phaseIn > 180) ? maxVal : minVal;
            end
        end
    endfunction

    always_ff @(posedge clock or posedge reset) begin
        if (reset || phase != prev_phase) begin
            tableSize <= logic_table_size; // Assign constant table size on reset
            prev_phase <= phase; // Update previous phase

            // Convert input phase into table index
            phaseIdx = phase_to_phaseVal(phase);
            phaseIdxOut <= phaseIdx;
            // Set initial index based on phase offset
            i <= calculate_start_index(phaseIdx);

            // Set initial traversal direction based on phase value
            if (phase >= 0) begin
                case (phase)
                    90: begin
                        // At 90º, reverse traversal
                        reverseTraversal <= 1;
                    end
                    180: begin
                        // At 180º, reverse traversal
                        reverseTraversal <= 1;
                    end
                    default: begin
                        // General case: forward traversal
                        reverseTraversal <= (i < `TABLE_SIZE - 1) ? 0 : 1;
                    end
                endcase
            end else begin
                case (phase)
                    -90: begin
                        // At -90º, forward traversal
                        reverseTraversal <= 0;
                    end
                    -180: begin
                        // At -180º, reverse traversal
                        reverseTraversal <= 1;
                    end
                    default: begin
                        // General case: reverse traversal
                        reverseTraversal <= (i > 0) ? 1 : 0;
                    end
                endcase
            end

            sine <= sine_wave_table[i]; // Initial output

        end else begin
            // Output current sine wave sample
            sine <= sine_wave_table[i];

            // Update index based on traversal direction
            if (!reverseTraversal) begin // Forward traversal
                if (i == tableSize - 1) begin
                    reverseTraversal <= 1; // Switch to reverse traversal at the end
                end 
                i <= i + 1; // Continue moving forward
            end else begin // Reverse traversal
                if (i == 1) begin
                    reverseTraversal <= 0; // Switch to forward traversal at the start
                end
                i <= i - 1; // Continue moving back
            end
        end
    end
endmodule
